library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

use work.top_level_types.all;


entity block_ram_4k is
	port(
		clk_0: in std_logic;
		port_0: in bram_port_32b;
		p0_read_data: out std_logic_vector(31 downto 0);
		
		clk_1: in std_logic;
		port_1: in bram_port_32b;
		p1_read_data: out std_logic_vector(31 downto 0)
	);
end block_ram_4k;

architecture Behavioral of block_ram_4k is
	signal p0_bram_address: std_logic_vector(13 downto 0) := (others => '0');
	signal p0_write_mask_0: std_logic_vector(0 to 3) := "0000";
	signal p0_write_mask_1: std_logic_vector(0 to 3) := "0000";
	signal p0_bram_select: std_logic_vector(0 downto 0) := "0";

	signal p0_data_out_0: std_logic_vector(31 downto 0) := (others => '0');
	signal p0_data_out_1: std_logic_vector(31 downto 0) := (others => '0');

	signal p1_bram_address: std_logic_vector(13 downto 0) := (others => '0');
	signal p1_write_mask_0: std_logic_vector(0 to 3) := "0000";
	signal p1_write_mask_1: std_logic_vector(0 to 3) := "0000";
	signal p1_bram_select: std_logic_vector(0 downto 0) := "0";

	signal p1_data_out_0: std_logic_vector(31 downto 0) := (others => '0');
	signal p1_data_out_1: std_logic_vector(31 downto 0) := (others => '0');

begin
	p0_bram_address <= port_0.address(10 downto 2) & "00000";
	p0_write_mask_0 <= port_0.write_mask when port_0.address(11) = '0' else "0000";
	p0_write_mask_1 <= port_0.write_mask when port_0.address(11) = '1' else "0000";
	p0_read_data <= p0_data_out_0 when p0_bram_select = "0" else p0_data_out_1;

	p1_bram_address <= port_1.address(10 downto 2) & "00000";
	p1_write_mask_0 <= port_1.write_mask when port_1.address(11) = '0' else "0000";
	p1_write_mask_1 <= port_1.write_mask when port_1.address(11) = '1' else "0000";
	p1_read_data <= p1_data_out_0 when p1_bram_select = "0" else p1_data_out_1;

	bram0 : RAMB16BWER
	generic map (
		-- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
		DATA_WIDTH_A => 36,
		DATA_WIDTH_B => 36,
		-- DOA_REG/DOB_REG: Optional output register (0 or 1)
		DOA_REG => 0,
		DOB_REG => 0,
		-- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
		EN_RSTRAM_A => FALSE,
		EN_RSTRAM_B => FALSE,
		-- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- INIT_A/INIT_B: Initial values on output port
		INIT_A => X"000000000",
		INIT_B => X"000000000",
		-- INIT_FILE: Optional file used to specify initial RAM contents
		INIT_FILE => "NONE",
		-- RSTTYPE: "SYNC" or "ASYNC"
		RSTTYPE => "SYNC",
		-- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR"
		RST_PRIORITY_A => "CE",
		RST_PRIORITY_B => "CE",
		-- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
		SIM_COLLISION_CHECK => "ALL",
		-- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
		SIM_DEVICE => "SPARTAN6",
		-- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
		SRVAL_A => X"000000000",
		SRVAL_B => X"000000000",
		-- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
		WRITE_MODE_A => "READ_FIRST",
		WRITE_MODE_B => "READ_FIRST"
	)
	port map (
		-- Port A Data: 32-bit (each) output: Port A data
		DOA => p0_data_out_0, -- 32-bit output: A port data output
		DOPA => open, -- 4-bit output: A port parity output
		-- Port B Data: 32-bit (each) output: Port B data
		DOB => p1_data_out_0, -- 32-bit output: B port data output
		DOPB => open, -- 4-bit output: B port parity output

		-- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
		ADDRA => p0_bram_address, -- 14-bit input: A port address input
		CLKA => clk_0, -- 1-bit input: A port clock input
		ENA => '1', -- 1-bit input: A port enable input
		REGCEA => '1', -- 1-bit input: A port register clock enable input
		RSTA => '0', -- 1-bit input: A port register set/reset input
		WEA => p0_write_mask_0, -- 4-bit input: Port A byte-wide write enable input
		-- Port A Data: 32-bit (each) input: Port A data
		DIA => port_0.write_data, -- 32-bit input: A port data input
		DIPA => (others => '0'), -- 4-bit input: A port parity input

		-- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
		ADDRB => p1_bram_address, -- 14-bit input: B port address input
		CLKB => clk_1, -- 1-bit input: B port clock input
		ENB => '1', -- 1-bit input: B port enable input
		REGCEB => '1', -- 1-bit input: B port register clock enable input
		RSTB => '0', -- 1-bit input: B port register set/reset input
		WEB => p1_write_mask_0, -- 4-bit input: Port B byte-wide write enable input
		-- Port B Data: 32-bit (each) input: Port B data
		DIB => port_1.write_data, -- 32-bit input: B port data input
		DIPB => (others => '0') -- 4-bit input: B port parity input
	);

	bram1 : RAMB16BWER
	generic map (
		-- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
		DATA_WIDTH_A => 36,
		DATA_WIDTH_B => 36,
		-- DOA_REG/DOB_REG: Optional output register (0 or 1)
		DOA_REG => 0,
		DOB_REG => 0,
		-- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
		EN_RSTRAM_A => FALSE,
		EN_RSTRAM_B => FALSE,
		-- INITP_00 to INITP_07: Initial memory contents.
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- INIT_00 to INIT_3F: Initial memory contents.
		INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- INIT_A/INIT_B: Initial values on output port
		INIT_A => X"000000000",
		INIT_B => X"000000000",
		-- INIT_FILE: Optional file used to specify initial RAM contents
		INIT_FILE => "NONE",
		-- RSTTYPE: "SYNC" or "ASYNC"
		RSTTYPE => "SYNC",
		-- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR"
		RST_PRIORITY_A => "CE",
		RST_PRIORITY_B => "CE",
		-- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
		SIM_COLLISION_CHECK => "ALL",
		-- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
		SIM_DEVICE => "SPARTAN6",
		-- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
		SRVAL_A => X"000000000",
		SRVAL_B => X"000000000",
		-- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
		WRITE_MODE_A => "READ_FIRST",
		WRITE_MODE_B => "READ_FIRST"
	)
	port map (
		-- Port A Data: 32-bit (each) output: Port A data
		DOA => p0_data_out_1, -- 32-bit output: A port data output
		DOPA => open, -- 4-bit output: A port parity output
		-- Port B Data: 32-bit (each) output: Port B data
		DOB => p1_data_out_1, -- 32-bit output: B port data output
		DOPB => open, -- 4-bit output: B port parity output

		-- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
		ADDRA => p0_bram_address, -- 14-bit input: A port address input
		CLKA => clk_0, -- 1-bit input: A port clock input
		ENA => '1', -- 1-bit input: A port enable input
		REGCEA => '1', -- 1-bit input: A port register clock enable input
		RSTA => '0', -- 1-bit input: A port register set/reset input
		WEA => p0_write_mask_1, -- 4-bit input: Port A byte-wide write enable input
		-- Port A Data: 32-bit (each) input: Port A data
		DIA => port_0.write_data, -- 32-bit input: A port data input
		DIPA => (others => '0'), -- 4-bit input: A port parity input

		-- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
		ADDRB => p1_bram_address, -- 14-bit input: B port address input
		CLKB => clk_1, -- 1-bit input: B port clock input
		ENB => '1', -- 1-bit input: B port enable input
		REGCEB => '1', -- 1-bit input: B port register clock enable input
		RSTB => '0', -- 1-bit input: B port register set/reset input
		WEB => p1_write_mask_1, -- 4-bit input: Port B byte-wide write enable input
		-- Port B Data: 32-bit (each) input: Port B data
		DIB => (port_1.write_data), -- 32-bit input: B port data input
		DIPB => (others => '0') -- 4-bit input: B port parity input
	);
	

	process(clk_0)
		variable v_opcode: std_logic_vector(31 downto 0);
	begin
		if rising_edge(clk_0) then
			p0_bram_select <= port_0.address(11 downto 11);
		end if;
	end process;

	process(clk_1)
		variable v_opcode: std_logic_vector(31 downto 0);
	begin
		if rising_edge(clk_1) then
			p1_bram_select <= port_1.address(11 downto 11);
		end if;
	end process;
end Behavioral;
