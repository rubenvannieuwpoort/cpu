library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.top_level_types.all;


entity textmode_vga_generator is
	port(
		clk: in std_logic;
		textbuffer_read_port_out: out bram_port_8b;
		textbuffer_read_data_in: in std_logic_vector(7 downto 0);
		--font_read_port_out: out bram_port_8b;
		--font_read_data_in: in std_logic_vector(7 downto 0);
		vga_out: out vga_signals
	);
end textmode_vga_generator;

-- VGA timings for different resolutions

-- HDTV (1280x720@60)
-- pixel clock: 74.2 MHz
-- 1280 72 80 216, 720 3 5 22

-- SDTV (720x480@60)
-- pixel clock: 27.7 MHz
-- 720 24 40 96, 480 10 3 32

-- VGA (640x480@60)
-- pixel clock: 27.17
-- 640 16 96 48, 480 10 2 33

architecture Behavioral of textmode_vga_generator is

	-- change this block to change the resolution
	-- you also need to change the frequency of the pixel clock
	constant width: natural := 1280;
	constant hFrontPorch: natural := 72;
	constant hSync: natural := 80;
	constant hBackPorch: natural := 216;

	constant height: natural := 720;
	constant vFrontPorch: natural := 3;
	constant vSync: natural := 5;
	constant vBackPorch: natural := 22;
	-- don't touch stuff after this line

	constant hSyncStart: natural := width + hFrontPorch;
	constant hSyncEnd: natural := hSyncStart + hSync;
	constant hMax: natural := hSyncEnd + hBackPorch - 1;
	constant hSyncActive: std_logic := '1';
	constant vSyncStart: natural := height + vFrontPorch;
	constant vSyncEnd: natural := vSyncStart + vSync;
	constant vMax: natural := vSyncEnd + vBackPorch - 1;
	
	constant characters_per_row: natural := 160;

	signal p: std_logic := '0';
	signal char_idx: unsigned(12 downto 0) := (others => '0');
	signal char_idx_base: unsigned(12 downto 0) := (others => '0');
	signal char: unsigned(7 downto 0) := (others => '0');
	signal x, x_1, x_2, x_3, x_4: unsigned(10 downto 0) := (others => '0');
	signal y, y_1, y_2, y_3, y_4: unsigned(10 downto 0) := (others => '0');

	type character_data is array(0 to 4095) of std_logic_vector(7 downto 0);

	constant font_data: character_data := (
	   -- Code page 437
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	   "00000000", "00000000", "01111110", "10000001", "10100101", "10000001", "10000001", "10111101", "10011001", "10000001", "10000001", "01111110", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "01111110", "11111111", "11011011", "11111111", "11111111", "11000011", "11100111", "11111111", "11111111", "01111110", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00110110", "01111111", "01111111", "01111111", "01111111", "00111110", "00011100", "00001000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00001000", "00011100", "00111110", "01111111", "00111110", "00011100", "00001000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00011000", "00111100", "00111100", "11100111", "11100111", "11100111", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00011000", "00111100", "01111110", "11111111", "11111111", "01111110", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011000", "00111100", "00111100", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11100111", "11000011", "11000011", "11100111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111100", "01100110", "01000010", "01000010", "01100110", "00111100", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "11111111", "11111111", "11111111", "11111111", "11111111", "11000011", "10011001", "10111101", "10111101", "10011001", "11000011", "11111111", "11111111", "11111111", "11111111", "11111111", -- ?
	   "00000000", "00000000", "01111000", "01110000", "01011000", "01001100", "00011110", "00110011", "00110011", "00110011", "00110011", "00011110", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00111100", "01100110", "01100110", "01100110", "00111100", "00011000", "01111110", "00011000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "11111100", "11001100", "11111100", "00001100", "00001100", "00001100", "00001100", "00001110", "00001111", "00000111", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "11111110", "11000110", "11111110", "11000110", "11000110", "11000110", "11000110", "11100110", "11100111", "01100111", "00000011", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00011000", "11011011", "01111110", "00111100", "01100110", "01100110", "00111100", "01111110", "11011011", "00011000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000001", "00000011", "00000111", "00001111", "00011111", "01111111", "00011111", "00001111", "00000111", "00000011", "00000001", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "01000000", "01100000", "01110000", "01111000", "01111100", "01111111", "01111100", "01111000", "01110000", "01100000", "01000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00011000", "00111100", "01111110", "00011000", "00011000", "00011000", "00011000", "01111110", "00111100", "00011000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "00000000", "01100110", "01100110", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "11111110", "11011011", "11011011", "11011011", "11011110", "11011000", "11011000", "11011000", "11011000", "11011000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00111110", "01100011", "00000110", "00011100", "00110110", "01100011", "01100011", "00110110", "00011100", "00110000", "01100011", "00111110", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "01111111", "01111111", "01111111", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00011000", "00111100", "01111110", "00011000", "00011000", "00011000", "01111110", "00111100", "00011000", "01111110", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00011000", "00111100", "01111110", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "01111110", "00111100", "00011000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00011000", "00110000", "01111111", "00110000", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00001100", "00000110", "01111111", "00000110", "00001100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000011", "00000011", "00000011", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00100100", "01100110", "11111111", "01100110", "00100100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00001000", "00011100", "00011100", "00111110", "00111110", "01111111", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "01111111", "01111111", "00111110", "00111110", "00011100", "00011100", "00001000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", --  
	   "00000000", "00000000", "00011000", "00111100", "00111100", "00111100", "00111100", "00011000", "00011000", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- !
	   "00000000", "01100110", "01100110", "01100110", "00100100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- "
	   "00000000", "00000000", "00110110", "00110110", "00110110", "01111111", "00110110", "00110110", "01111111", "00110110", "00110110", "00110110", "00000000", "00000000", "00000000", "00000000", -- #
	   "00011000", "00011000", "00111110", "01100011", "01000011", "00000011", "00111110", "01100000", "01100000", "01100001", "01100011", "00111110", "00011000", "00011000", "00000000", "00000000", -- $
	   "00000000", "00000000", "00000000", "00000000", "01000011", "01100011", "00110000", "00011000", "00001100", "00000110", "01100011", "01100001", "00000000", "00000000", "00000000", "00000000", -- %
	   "00000000", "00000000", "00011100", "00110110", "00110110", "00011100", "01101110", "00111011", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- &&
	   "00000000", "00001100", "00001100", "00001100", "00000110", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- '
	   "00000000", "00000000", "00110000", "00011000", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00011000", "00110000", "00000000", "00000000", "00000000", "00000000", -- (
	   "00000000", "00000000", "00001100", "00011000", "00110000", "00110000", "00110000", "00110000", "00110000", "00110000", "00011000", "00001100", "00000000", "00000000", "00000000", "00000000", -- )
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01100110", "00111100", "11111111", "00111100", "01100110", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- *
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "01111110", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "00011000", "00001100", "00000000", "00000000", "00000000", -- ,
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- -
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- .
	   "00000000", "00000000", "00000000", "00000000", "01000000", "01100000", "00110000", "00011000", "00001100", "00000110", "00000011", "00000001", "00000000", "00000000", "00000000", "00000000", -- /
	   "00000000", "00000000", "01111110", "11000011", "11000011", "11000011", "11011011", "11011011", "11000011", "11000011", "11000011", "01111110", "00000000", "00000000", "00000000", "00000000", -- 0
	   "00000000", "00000000", "00011000", "00011110", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "01111110", "00000000", "00000000", "00000000", "00000000", -- 1
	   "00000000", "00000000", "00111110", "01100011", "01100011", "01100000", "00110000", "00011000", "00001100", "00000110", "01100011", "01111111", "00000000", "00000000", "00000000", "00000000", -- 2
	   "00000000", "00000000", "00111110", "01100011", "01100000", "01100000", "00111100", "01100000", "01100000", "01100000", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- 3
	   "00000000", "00000000", "00110000", "00111000", "00111100", "00110110", "00110011", "00110011", "01111111", "00110000", "00110000", "01111000", "00000000", "00000000", "00000000", "00000000", -- 4
	   "00000000", "00000000", "01111111", "00000011", "00000011", "00000011", "00111111", "01100000", "01100000", "01100000", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- 5
	   "00000000", "00000000", "00111110", "00000011", "00000011", "00000011", "00111111", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- 6
	   "00000000", "00000000", "01111111", "01100011", "01100000", "00110000", "00011000", "00001100", "00001100", "00001100", "00001100", "00001100", "00000000", "00000000", "00000000", "00000000", -- 7
	   "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "00111110", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- 8
	   "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01111110", "01100000", "01100000", "01100000", "00111110", "00000000", "00000000", "00000000", "00000000", -- 9
	   "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", -- :
	   "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00011000", "00011000", "00001100", "00000000", "00000000", "00000000", "00000000", -- ;
	   "00000000", "00000000", "00000000", "01100000", "00110000", "00011000", "00001100", "00000110", "00001100", "00011000", "00110000", "01100000", "00000000", "00000000", "00000000", "00000000", -- <
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "00000000", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- =
	   "00000000", "00000000", "00000000", "00000110", "00001100", "00011000", "00110000", "01100000", "00110000", "00011000", "00001100", "00000110", "00000000", "00000000", "00000000", "00000000", -- >
	   "00000000", "00000000", "00111110", "01100011", "01100011", "00110000", "00011000", "00011000", "00011000", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- ?
	   "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01111011", "01111011", "01111011", "00111011", "00000011", "01111110", "00000000", "00000000", "00000000", "00000000", -- @
	   "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01111111", "01100011", "01100011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- A
	   "00000000", "00000000", "00111111", "01100110", "01100110", "01100110", "00111110", "01100110", "01100110", "01100110", "01100110", "00111111", "00000000", "00000000", "00000000", "00000000", -- B
	   "00000000", "00000000", "00111110", "01100011", "01000011", "00000011", "00000011", "00000011", "00000011", "01000011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- C
	   "00000000", "00000000", "00111111", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "00111111", "00000000", "00000000", "00000000", "00000000", -- D
	   "00000000", "00000000", "01111111", "01100110", "00000110", "00100110", "00111110", "00100110", "00000110", "00000110", "01100110", "01111111", "00000000", "00000000", "00000000", "00000000", -- E
	   "00000000", "00000000", "01111111", "01100110", "00000110", "00100110", "00111110", "00100110", "00000110", "00000110", "00000110", "00001111", "00000000", "00000000", "00000000", "00000000", -- F
	   "00000000", "00000000", "00111110", "01100011", "01100011", "00000011", "00000011", "01111011", "01100011", "01100011", "01100011", "01011110", "00000000", "00000000", "00000000", "00000000", -- G
	   "00000000", "00000000", "01100011", "01100011", "01100011", "01100011", "01111111", "01100011", "01100011", "01100011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- H
	   "00000000", "00000000", "01111110", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "01111110", "00000000", "00000000", "00000000", "00000000", -- I
	   "00000000", "00000000", "01111000", "00110000", "00110000", "00110000", "00110000", "00110000", "00110011", "00110011", "00110011", "00011110", "00000000", "00000000", "00000000", "00000000", -- J
	   "00000000", "00000000", "01100011", "01100011", "00110011", "00011011", "00001111", "00001111", "00011011", "00110011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- K
	   "00000000", "00000000", "00001111", "00000110", "00000110", "00000110", "00000110", "00000110", "00000110", "01000110", "01100110", "01111111", "00000000", "00000000", "00000000", "00000000", -- L
	   "00000000", "00000000", "11000011", "11100111", "11111111", "11111111", "11011011", "11000011", "11000011", "11000011", "11000011", "11000011", "00000000", "00000000", "00000000", "00000000", -- M
	   "00000000", "00000000", "01100011", "01100011", "01100111", "01100111", "01101111", "01111011", "01110011", "01110011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- N
	   "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- O
	   "00000000", "00000000", "00111111", "01100110", "01100110", "01100110", "01100110", "00111110", "00000110", "00000110", "00000110", "00001111", "00000000", "00000000", "00000000", "00000000", -- P
	   "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01101011", "01111011", "00111110", "00110000", "01110000", "00000000", "00000000", -- Q
	   "00000000", "00000000", "00111111", "01100110", "01100110", "01100110", "00111110", "00110110", "01100110", "01100110", "01100110", "01100111", "00000000", "00000000", "00000000", "00000000", -- R
	   "00000000", "00000000", "00111110", "01100011", "00000011", "00000011", "00001110", "00111000", "01100000", "01100000", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- S
	   "00000000", "00000000", "11111111", "11011011", "10011001", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- T
	   "00000000", "00000000", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- U
	   "00000000", "00000000", "11000011", "11000011", "11000011", "11000011", "11000011", "11000011", "11000011", "01100110", "00111100", "00011000", "00000000", "00000000", "00000000", "00000000", -- V
	   "00000000", "00000000", "11000011", "11000011", "11000011", "11000011", "11000011", "11011011", "11011011", "11111111", "11100111", "11000011", "00000000", "00000000", "00000000", "00000000", -- W
	   "00000000", "00000000", "11000011", "11000011", "11000011", "01100110", "00111100", "00111100", "01100110", "11000011", "11000011", "11000011", "00000000", "00000000", "00000000", "00000000", -- X
	   "00000000", "00000000", "11000011", "11000011", "11000011", "11000011", "01100110", "00111100", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- Y
	   "00000000", "00000000", "01111111", "01100011", "01100001", "00110000", "00011000", "00001100", "00000110", "01000011", "01100011", "01111111", "00000000", "00000000", "00000000", "00000000", -- Z
	   "00000000", "00000000", "00111100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00001100", "00111100", "00000000", "00000000", "00000000", "00000000", -- p
	   "00000000", "00000000", "00000000", "00000001", "00000011", "00000111", "00001110", "00011100", "00111000", "01110000", "01100000", "01000000", "00000000", "00000000", "00000000", "00000000", -- \
	   "00000000", "00000000", "00111100", "00110000", "00110000", "00110000", "00110000", "00110000", "00110000", "00110000", "00110000", "00111100", "00000000", "00000000", "00000000", "00000000", -- ]
	   "00000000", "00001000", "00011100", "00110110", "01100011", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ^
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "00000000", "00000000", -- _
	   "00000000", "00001100", "00001100", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- `
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00011110", "00110000", "00111110", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- a
	   "00000000", "00000000", "00000111", "00000110", "00000110", "00111110", "01100110", "01100110", "01100110", "01100110", "01100110", "00111111", "00000000", "00000000", "00000000", "00000000", -- b
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111110", "01100011", "00000011", "00000011", "00000011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- c
	   "00000000", "00000000", "00111000", "00110000", "00110000", "00111110", "00110011", "00110011", "00110011", "00110011", "00110011", "01111110", "00000000", "00000000", "00000000", "00000000", -- d
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111110", "01100011", "01100011", "01111111", "00000011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- e
	   "00000000", "00000000", "00111000", "01101100", "00001100", "00001100", "00111111", "00001100", "00001100", "00001100", "00001100", "00011110", "00000000", "00000000", "00000000", "00000000", -- f
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01101110", "00110011", "00110011", "00110011", "00110011", "00110011", "00111110", "00110000", "00110011", "00011110", "00000000", -- g
	   "00000000", "00000000", "00000111", "00000110", "00000110", "00111110", "01100110", "01100110", "01100110", "01100110", "01100110", "01100111", "00000000", "00000000", "00000000", "00000000", -- h
	   "00000000", "00000000", "00011000", "00011000", "00000000", "00011100", "00011000", "00011000", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- i
	   "00000000", "00000000", "00110000", "00110000", "00000000", "00111000", "00110000", "00110000", "00110000", "00110000", "00110000", "00110000", "00110011", "00110011", "00011110", "00000000", -- j
	   "00000000", "00000000", "00000111", "00000110", "00000110", "01100110", "00110110", "00011110", "00011110", "00110110", "01100110", "01100111", "00000000", "00000000", "00000000", "00000000", -- k
	   "00000000", "00000000", "00011100", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- l
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01100111", "11111111", "11011011", "11011011", "11011011", "11000011", "11000011", "00000000", "00000000", "00000000", "00000000", -- m
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111011", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "00000000", "00000000", "00000000", "00000000", -- n
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- o
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111011", "01100110", "01100110", "01100110", "01100110", "01100110", "00111110", "00000110", "00000110", "00001111", "00000000", -- p
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01101110", "00110011", "00110011", "00110011", "00110011", "00110011", "00111110", "00110000", "00110000", "01111000", "00000000", -- q
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111011", "01101110", "01100110", "00000110", "00000110", "00000110", "00001111", "00000000", "00000000", "00000000", "00000000", -- r
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00111110", "01100011", "00000011", "00111110", "01100000", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- s
	   "00000000", "00000000", "00001100", "00001100", "00001100", "00111111", "00001100", "00001100", "00001100", "00001100", "01101100", "00111000", "00000000", "00000000", "00000000", "00000000", -- t
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00110011", "00110011", "00110011", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- u
	   "00000000", "00000000", "00000000", "00000000", "00000000", "11000011", "11000011", "11000011", "11000011", "01100110", "00111100", "00011000", "00000000", "00000000", "00000000", "00000000", -- v
	   "00000000", "00000000", "00000000", "00000000", "00000000", "11000011", "11000011", "11011011", "11011011", "11011011", "11111111", "01100110", "00000000", "00000000", "00000000", "00000000", -- w
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01100011", "01100011", "00110110", "00011100", "00110110", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- x
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01111110", "01100000", "00110000", "00011111", "00000000", -- y
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "01100001", "00110000", "00011000", "00001100", "01000110", "01111111", "00000000", "00000000", "00000000", "00000000", -- z
	   "00000000", "00000000", "01110000", "00011000", "00011000", "00011000", "00001110", "00011000", "00011000", "00011000", "00011000", "01110000", "00000000", "00000000", "00000000", "00000000", -- {
	   "00000000", "00000000", "00011000", "00011000", "00011000", "00011000", "00000000", "00011000", "00011000", "00011000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- |
	   "00000000", "00000000", "00001110", "00011000", "00011000", "00011000", "01110000", "00011000", "00011000", "00011000", "00011000", "00001110", "00000000", "00000000", "00000000", "00000000", -- }
	   "00000000", "00000000", "01101110", "00111011", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- ~
	   "00000000", "00000000", "00000000", "00000000", "00001000", "00011100", "00110110", "01100011", "01100011", "01100011", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00111100", "01100110", "01000011", "00000011", "00000011", "00000011", "01000011", "01100110", "00111100", "00110000", "01100000", "00111110", "00000000", "00000000", -- �
	   "00000000", "00000000", "00110011", "00000000", "00000000", "00110011", "00110011", "00110011", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00110000", "00011000", "00001100", "00000000", "00111110", "01100011", "01100011", "01111111", "00000011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00001100", "00011110", "00110011", "00000000", "00011110", "00110000", "00111110", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00110011", "00000000", "00000000", "00011110", "00110000", "00111110", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000110", "00001100", "00011000", "00000000", "00011110", "00110000", "00111110", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00011100", "00110110", "00011100", "00000000", "00011110", "00110000", "00111110", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00111110", "01100011", "00000011", "00000011", "01100011", "00111110", "00011000", "00110000", "00110110", "00011100", "00000000", "00000000", -- �
	   "00000000", "00001100", "00011110", "00110011", "00000000", "00111110", "01100011", "01100011", "01111111", "00000011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00110011", "00000000", "00000000", "00111110", "01100011", "01100011", "01111111", "00000011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000110", "00001100", "00011000", "00000000", "00111110", "01100011", "01100011", "01111111", "00000011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "01100110", "00000000", "00000000", "00011100", "00011000", "00011000", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00011000", "00111100", "01100110", "00000000", "00011100", "00011000", "00011000", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000110", "00001100", "00011000", "00000000", "00011100", "00011000", "00011000", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "01100011", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01111111", "01100011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- �
	   "00011100", "00110110", "00011100", "00000000", "00111110", "01100011", "01100011", "01100011", "01111111", "01100011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- �
	   "00110000", "00011000", "00001100", "00000000", "01111111", "01100110", "00000110", "00111110", "00000110", "00000110", "01100110", "01111111", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "01100110", "11011011", "11011000", "11111110", "00011011", "00011011", "11111011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "01111110", "00011011", "00011011", "00011011", "00011011", "01111111", "00011011", "00011011", "00011011", "01111011", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00001100", "00011110", "00110011", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "01100011", "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000110", "00001100", "00011000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00001100", "00011110", "00110011", "00000000", "00110011", "00110011", "00110011", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000110", "00001100", "00011000", "00000000", "00110011", "00110011", "00110011", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "01100011", "00000000", "00000000", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01111110", "01100000", "00110000", "00011111", "00000000", -- �
	   "00000000", "01100011", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "01100011", "00000000", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00011000", "00011000", "00111110", "01100011", "00000011", "00000011", "01100011", "00111110", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00011100", "00110110", "00100110", "00000110", "00001111", "00000110", "00000110", "00000110", "00000110", "01100111", "00111111", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "11000011", "01100110", "00111100", "00011000", "11111111", "00011000", "11111111", "00011000", "00011000", "00011000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00111111", "01100011", "01100011", "00111111", "00000011", "00110011", "01111011", "00110011", "00110011", "00110011", "01100011", "00000000", "00000000", "00000000", "00000000", -- P
	   "00000000", "01110000", "11011000", "00011000", "00011000", "00011000", "01111110", "00011000", "00011000", "00011000", "00011000", "00011000", "00011011", "00001110", "00000000", "00000000", -- �
	   "00000000", "00110000", "00011000", "00001100", "00000000", "00011110", "00110000", "00111110", "00110011", "00110011", "00111011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00110000", "00011000", "00001100", "00000000", "00011100", "00011000", "00011000", "00011000", "00011000", "00011000", "00111100", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00110000", "00011000", "00001100", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00011000", "00001100", "00000110", "00000000", "00110011", "00110011", "00110011", "00110011", "00110011", "00110011", "01101110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "01101110", "00111011", "00000000", "00111011", "01100110", "01100110", "01100110", "01100110", "01100110", "01100110", "00000000", "00000000", "00000000", "00000000", -- �
	   "01101110", "00111011", "00000000", "01100011", "01100111", "01101111", "01111111", "01111011", "01110011", "01100011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00111100", "00110110", "00110110", "01111100", "00000000", "01111110", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00011100", "00110110", "00110110", "00011100", "00000000", "00111110", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00001100", "00001100", "00000000", "00001100", "00001100", "00001100", "00000110", "01100011", "01100011", "00111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "00000011", "00000011", "00000011", "00000011", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "01100000", "01100000", "01100000", "01100000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000110", "00000110", "01000110", "01100110", "00110110", "00011000", "00001100", "00000110", "00111011", "01101101", "00110000", "00011000", "01111100", "00000000", "00000000", -- �
	   "00000000", "00000110", "00000110", "01000110", "01100110", "00110110", "00011000", "00001100", "01100110", "01110011", "01101001", "01111100", "01100000", "01100000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00011000", "00011000", "00000000", "00011000", "00011000", "00111100", "00111100", "00111100", "00111100", "00011000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01101100", "00110110", "00011011", "00110110", "01101100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00011011", "00110110", "01101100", "00110110", "00011011", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "10001000", "00100010", "10001000", "00100010", "10001000", "00100010", "10001000", "00100010", "10001000", "00100010", "10001000", "00100010", "10001000", "00100010", "10001000", "00100010", -- �
	   "01010101", "10101010", "01010101", "10101010", "01010101", "10101010", "01010101", "10101010", "01010101", "10101010", "01010101", "10101010", "01010101", "10101010", "01010101", "10101010", -- �
	   "10111011", "11101110", "10111011", "11101110", "10111011", "11101110", "10111011", "11101110", "10111011", "11101110", "10111011", "11101110", "10111011", "11101110", "10111011", "11101110", -- �
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- �
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- �
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011111", "00011000", "00011111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- �
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011000", "00011111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- +
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101111", "01100000", "01101111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- �
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01111111", "01100000", "01101111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- +
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101111", "01100000", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011111", "00011000", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "11111000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- -
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- -
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "11111000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- -
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "11111111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "11111000", "00011000", "11111000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- �
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "11101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- �
	   "01101100", "01101100", "01101100", "01101100", "01101100", "11101100", "00001100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00001100", "11101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- +
	   "01101100", "01101100", "01101100", "01101100", "01101100", "11101111", "00000000", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- -
	   "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "00000000", "11101111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- -
	   "01101100", "01101100", "01101100", "01101100", "01101100", "11101100", "00001100", "11101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "00000000", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- -
	   "01101100", "01101100", "01101100", "01101100", "01101100", "11101111", "00000000", "11101111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "11111111", "00000000", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- -
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- -
	   "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "00000000", "11111111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- -
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- -
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "11111000", "00011000", "11111000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "11111000", "00011000", "11111000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- +
	   "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "11111111", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", "01101100", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "11111111", "00011000", "11111111", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- +
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- +
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- +
	   "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", -- _
	   "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", "00001111", -- �
	   "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", "11110000", -- �
	   "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01101110", "00111011", "00011011", "00011011", "00011011", "00111011", "01101110", "00000000", "00000000", "00000000", "00000000", -- a
	   "00000000", "00000000", "00011110", "00110011", "00110011", "00110011", "00011011", "00110011", "01100011", "01100011", "01100011", "00110011", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "01111111", "01100011", "01100011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000011", "00000000", "00000000", "00000000", "00000000", -- G
	   "00000000", "00000000", "00000000", "00000000", "01111111", "00110110", "00110110", "00110110", "00110110", "00110110", "00110110", "00110110", "00000000", "00000000", "00000000", "00000000", -- p
	   "00000000", "00000000", "00000000", "01111111", "01100011", "00000110", "00001100", "00011000", "00001100", "00000110", "01100011", "01111111", "00000000", "00000000", "00000000", "00000000", -- S
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01111110", "00011011", "00011011", "00011011", "00011011", "00011011", "00001110", "00000000", "00000000", "00000000", "00000000", -- s
	   "00000000", "00000000", "00000000", "00000000", "01100110", "01100110", "01100110", "01100110", "01100110", "00111110", "00000110", "00000110", "00000011", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "01101110", "00111011", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", -- t
	   "00000000", "00000000", "00000000", "01111110", "00011000", "00111100", "01100110", "01100110", "01100110", "00111100", "00011000", "01111110", "00000000", "00000000", "00000000", "00000000", -- F
	   "00000000", "00000000", "00000000", "00011100", "00110110", "01100011", "01100011", "01111111", "01100011", "01100011", "00110110", "00011100", "00000000", "00000000", "00000000", "00000000", -- T
	   "00000000", "00000000", "00011100", "00110110", "01100011", "01100011", "01100011", "00110110", "00110110", "00110110", "00110110", "01110111", "00000000", "00000000", "00000000", "00000000", -- O
	   "00000000", "00000000", "01111000", "00001100", "00011000", "00110000", "01111100", "01100110", "01100110", "01100110", "01100110", "00111100", "00000000", "00000000", "00000000", "00000000", -- d
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01111110", "11011011", "11011011", "11011011", "01111110", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- 8
	   "00000000", "00000000", "00000000", "11000000", "01100000", "01111110", "11011011", "11011011", "11001111", "01111110", "00000110", "00000011", "00000000", "00000000", "00000000", "00000000", -- f
	   "00000000", "00000000", "00111000", "00001100", "00000110", "00000110", "00111110", "00000110", "00000110", "00000110", "00001100", "00111000", "00000000", "00000000", "00000000", "00000000", -- e
	   "00000000", "00000000", "00000000", "00111110", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "01100011", "00000000", "00000000", "00000000", "00000000", -- n
	   "00000000", "00000000", "00000000", "00000000", "01111111", "00000000", "00000000", "01111111", "00000000", "00000000", "01111111", "00000000", "00000000", "00000000", "00000000", "00000000", -- =
	   "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "01111110", "00011000", "00011000", "00000000", "00000000", "01111110", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00001100", "00011000", "00110000", "01100000", "00110000", "00011000", "00001100", "00000000", "01111110", "00000000", "00000000", "00000000", "00000000", -- =
	   "00000000", "00000000", "00000000", "00110000", "00011000", "00001100", "00000110", "00001100", "00011000", "00110000", "00000000", "01111110", "00000000", "00000000", "00000000", "00000000", -- =
	   "00000000", "00000000", "01110000", "11011000", "11011000", "11011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", -- (
	   "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011000", "00011011", "00011011", "00011011", "00001110", "00000000", "00000000", "00000000", "00000000", -- )
	   "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "00000000", "01111110", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01101110", "00111011", "00000000", "01101110", "00111011", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00011110", "00110011", "00110011", "00011110", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011000", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "11110000", "00110000", "00110000", "00110000", "00110000", "00110000", "00110111", "00110110", "00110110", "00111100", "00111000", "00000000", "00000000", "00000000", "00000000", -- v
	   "00000000", "00011011", "00110110", "00110110", "00110110", "00110110", "00110110", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- n
	   "00000000", "00001110", "00011011", "00011000", "00001100", "00000110", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "01111110", "01111110", "01111110", "01111110", "01111110", "01111110", "00000000", "00000000", "00000000", "00000000", "00000000", -- �
	   "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000"
	);

	--type text_buffer_data is array(0 to 7199) of std_logic_vector(7 downto 0);
	--constant text_buffer: text_buffer_data := (
	--	"01001000", "01100101", "01101100", "01101100", "01101111", "00101100", "00100000", "01110111", "01101111", "01110010", "01101100", "01100100", "00100001", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
	--	"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "01100010", "01111001", "01100101"
	--);

begin
	textbuffer_read_port_out.write_data <= (others => '0');
	textbuffer_read_port_out.write_mask <= (others => '0');
	textbuffer_read_port_out.address <= std_logic_vector(char_idx);
	--font_read_port_out.write_data <= (others => '0');
	--font_read_port_out.write_mask <= (others => '0');
	--font_read_port_out.address(12) <= '0';
	--font_read_port_out.address(11 downto 4) <= textbuffer_read_data_in(7 downto 0);
	--font_read_port_out.address(3 downto 0) <= std_logic_vector(y_2(3 downto 0));

	process(clk)
		variable idx: std_logic_vector(11 downto 0);
		variable row: std_logic_vector(7 downto 0);
	begin
		if rising_edge(clk) then
			if x < width and y < height then
				if p = '1' then
					vga_out.red <= "111";
					vga_out.green <= "111";
					vga_out.blue <= "11";
				else
					vga_out.red <= "000";
					vga_out.green <= "000";
					vga_out.blue <= "00";
				end if;
			else
				vga_out.red <= "000";
				vga_out.green <= "000";
				vga_out.blue <= "00";
			end if;

			-- track horizontal and vertical position and generate sync pulses
			if x_3 < hMax then
				x_3 <= x_3 + 1;
				
				if x_3(2 downto 0) = "111" then
					char_idx <= char_idx + 1;
				end if;
			else
				x_3 <= (others => '0');
				if y_3 < vMax then
					y_3 <= y_3 + 1;
					
					if y_3(3 downto 0) = "1111" then
						char_idx <= char_idx_base + characters_per_row;
						char_idx_base <= char_idx_base + characters_per_row;
					else
						char_idx <= char_idx_base;
					end if;
				else
					y_3 <= (others => '0');
					char_idx <= (others => '0');
					char_idx_base <= (others => '0');
				end if;
			end if;
			
			--x_3 <= x_4;
			--y_3 <= y_4;
			
			x_2 <= x_3;
			y_2 <= y_3;

			x_1 <= x_2;
			y_1 <= y_2;

			x <= x_1;
			y <= y_1;

			-- char_idx is the index in the text buffer to look up
			-- `char` lags one cycle behind `x` and `y`
			-- char <= unsigned(text_buffer(to_integer(char_idx)));
			char <= unsigned(textbuffer_read_data_in);

			-- index of the character, to look up the font data
			idx := std_logic_vector(char & y_1(3 downto 0));

			-- one row of font data
			-- `row` and `p` lag two cycles behind `x` and `y`
			row := font_data(to_integer(unsigned(idx)));

			-- store pixel value; '0' if background, '1' if foreground
			p <= row(to_integer(unsigned(x_1(2 downto 0))));

			if vSyncStart <= y and y < vSyncEnd then
				vga_out.vsync <= '1';
			else
				vga_out.vsync <= '0';
			end if;

			if hSyncStart <= x and x < hSyncEnd then
				vga_out.hsync <= '1';
			else
				vga_out.hsync <= '0';
			end if;
		end if;
	end process;
end Behavioral;
